----------------------------------------------------------------------------------
-- USE WORK.pkg_types.ALL;
----------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.pkg_constants.all;
----------------------------------------------------------------------------------
PACKAGE pkg_types IS
----------------------------------------------------------------------------------

  TYPE type_pwm_ref IS ARRAY(G_NCH-1 DOWNTO 0) OF STD_LOGIC_VECTOR(G_RES-1 DOWNTO 0);

----------------------------------------------------------------------------------
END;
----------------------------------------------------------------------------------
