----------------------------------------------------------------------------------
-- USE WORK.pkg_constants.ALL;
----------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
----------------------------------------------------------------------------------
PACKAGE pkg_constants IS
----------------------------------------------------------------------------------

  CONSTANT G_NCH        : POSITIVE := 8;
  CONSTANT G_RES        : POSITIVE := 8;

----------------------------------------------------------------------------------
end;
----------------------------------------------------------------------------------
